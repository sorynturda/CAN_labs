[aimspice]
[description]
204
stabilizator parametric cu dioda Zener
D1 1 2 Dioda
D4 3 2 Dioda
D2 0 1 Dioda
D3 0 3 Dioda
R 0 2 100
C 0 2 1m
D5 0 2 Zener
.Model Dioda D !tt=1e-9
.Model Zener D bv=6.8
Vin 1 3 sin (0 10 50 0 0)
[tran]
1e-9
50e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -1.35589E-29 8
1
v(2)
[end]
