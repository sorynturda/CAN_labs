[aimspice]
[description]
145
redresor dubla alternanta
D1 1 2 Dioda
D4 3 2 Dioda
D2 0 1 Dioda
D3 0 3 Dioda
R 2 0 100
.Model Dioda D tt=1e-9

Vin 1 3 sin (0 10 1k 0 0)
[tran]
1e-8
60e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
[end]
