[aimspice]
[description]
152
redresor cu filtru
D1 1 2 Dioda
D4 3 2 Dioda
D2 0 1 Dioda
D3 0 3 Dioda
R 0 2 100
C 0 2 3m
.Model Dioda D !tt=1e-9

Vin 1 3 dc 5 sin(0 8 50 0 0)
[tran]
1e-8
60e-3
X
X
0
[ana]
4 0
[end]
