[aimspice]
[description]
203
inversor cmos
V1 dd 0 dc 5
V2 ss 0 dc 0
V3 in 0 dc pulse (0 5 0 1e-10 1e-10 1e-6 2e-6)
C1 out 0 0.1p
MP out in dd dd MOS1
MN out in ss ss MOS

.Model MOS nmos vto 1.5
.Model MOS1 pmos vto -1.5

[dc]
1
V3
0
5
0.1
[ana]
1 2
0
1 1
1 1 -1 6
2
v3
v(out)
0
1 1
1 1 -1.2E-05 0
1
i(v1)
[end]
